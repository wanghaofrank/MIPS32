module Adder4(s,pp,gg,a,b,ci,z);
input [3:0] a;
input [3:0] b;
input ci;
output pp,gg,z;
output [3:0] s;
wire c1,c2,c3;
wire [3:0] p;
wire [3:0] g;
assign p=a^b;
assign g=a&b;
assign s=p^{c3,c2,c1,ci};
assign c1=g[0]|(p[0]&ci);
assign c2=g[1]|(p[1]&g[0])|(p[1]&p[0]&ci);
assign c3=g[2]|(p[2]&g[1])|(p[2]&p[1]&g[0])|(p[2]&p[1]&p[0]&ci);
assign pp=&p;
assign gg=g[3]|(p[3]&g[2])|(p[3]&p[2]&g[1])|(p[3]&p[2]&p[1]&g[0]);
assign z=&((({4{ci}}|{b[2]|b[1]|b[0],b[1]|b[0],b[0],1'b1})^b)^(~a));
endmodule

module Adder4_v(s,co,v,a,b,ci,z);
input [3:0] a;
input [3:0] b;
input ci;
output co,v,z;
output [3:0] s;
wire c1,c2,c3;
wire [3:0] p;
wire [3:0] g;
assign p=a^b;
assign g=a&b;
assign s=p^{c3,c2,c1,ci};
assign c1=g[0]|(p[0]&ci);
assign c2=g[1]|(p[1]&g[0])|(p[1]&p[0]&ci);
assign c3=g[2]|(p[2]&g[1])|(p[2]&p[1]&g[0])|(p[2]&p[1]&p[0]&ci);
assign co=g[3]|(p[3]&g[2])|(p[3]&p[2]&g[1])|(p[3]&p[2]&p[1]&g[0])|(p[3]&p[2]&p[1]&p[0]&ci);
assign v=c3^co;
assign z=&((({4{ci}}|{b[2]|b[1]|b[0],b[1]|b[0],b[0],1'b1})^b)^(~a));
endmodule

module Adder(s,co,a,b,ci,v,zero);
input [31:0] a;
input [31:0] b;
input ci;
output co,v,zero;
output [31:0] s;
wire c1,c2,c3,c4,c5,c6,c7,p1,p2,p3,p4,p5,p6,p7,g1,g2,g3,g4,g5,g6,g7;
wire [7:0] z;
wire [3:0] s0;
wire [3:0] s1;
wire [3:0] s2;
wire [3:0] s3;
wire [3:0] s4;
wire [3:0] s5;
wire [3:0] s6;
wire [3:0] s7;
assign c1=g1|(p1&ci);
assign c2=g2|(p2&g1)|(p2&p1&ci);
assign c3=g3|(p3&g2)|(p3&p2&g1)|(p3&p2&p1&ci);
assign c4=g4|(p4&g3)|(p4&p3&g2)|(p4&p3&p2&g1)|(p4&p3&p2&p1&ci);
assign c5=g5|(p5&g4)|(p5&p4&g3)|(p5&p4&p3&g2)|(p5&p4&p3&p2&g1)|(p5&p4&p3&p2&p1&ci);
assign c6=g6|(p6&g5)|(p6&p5&g4)|(p6&p5&p4&g3)|(p6&p5&p4&p3&g2)|(p6&p5&p4&p3&p2&g1)|(p6&p5&p4&p3&p2&p1&ci);
assign c7=g7|(p7&g6)|(p7&p6&g5)|(p7&p6&p5&g4)|(p7&p6&p5&p4&g3)|(p7&p6&p5&p4&p3&g2)|(p7&p6&p5&p4&p3&p2&g1)|(p7&p6&p5&p4&p3&p2&p1&ci);
Adder4 a0(s0,p1,g1,a[3:0],b[3:0],ci,z[0]);
Adder4 a1(s1,p2,g2,a[7:4],b[7:4],c1,z[1]);
Adder4 a2(s2,p3,g3,a[11:8],b[11:8],c2,z[2]);
Adder4 a3(s3,p4,g4,a[15:12],b[15:12],c3,z[3]);
Adder4 a4(s4,p5,g5,a[19:16],b[19:16],c4,z[4]);
Adder4 a5(s5,p6,g6,a[23:20],b[23:20],c5,z[5]);
Adder4 a6(s6,p7,g7,a[27:24],b[27:24],c6,z[6]);
Adder4_v a7(s7,co,v,a[31:28],b[31:28],c7,z[7]);
assign s={s7,s6,s5,s4,s3,s2,s1,s0};
assign zero=&z;
endmodule